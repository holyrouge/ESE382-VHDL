-----------------------------------------------------------------------
--
-- Title       : programmable_prescalar_tb
-- Design      : programmable_prescalar_tb
-- Authors     : Prangon Ghose (111623211), Albert Thomas (111386879)
-- Company     : Stony Brook University
-- Date		   : 04/10/2019
-- Lab Section : 01
-- Bench Number: 05
-- Lab Number  : 08
--
-----------------------------------------------------------------------
--
-- Description : programmable_prescalar_tb is a testbench for the
-- programmable_prescalar. It was generated by Active-HDL from simulation
-- data based on stimulators.
--
-- Inputs: None
-- Outputs: None			 
-----------------------------------------------------------------------

library ieee;
use ieee.NUMERIC_STD.all;
use ieee.std_logic_1164.all;

	-- Add your library and packages declaration here ...

entity programmable_prescalar_tb is
	-- Generic declarations of the tested unit
end programmable_prescalar_tb;

architecture testbench of programmable_prescalar_tb is
	-- Component declaration of the tested unit
	component programmable_prescalar
	port(
		clear : in STD_LOGIC;
		clk : in STD_LOGIC;
		cs : in STD_LOGIC_VECTOR(2 downto 0);
		clk_prescaled : out STD_LOGIC );
	end component;

	-- Stimulus signals - signals mapped to the input and inout ports of tested entity
	signal clear : STD_LOGIC;
	signal clk : STD_LOGIC;
	signal cs : STD_LOGIC_VECTOR(2 downto 0);
	-- Observed signals - signals mapped to the output ports of tested entity
	signal clk_prescaled : STD_LOGIC;

	-- Add your code here ...

begin

	-- Unit Under Test port map
	UUT : programmable_prescalar
		port map (
			clear => clear,
			clk => clk,
			cs => cs,
			clk_prescaled => clk_prescaled
		);

	--Below VHDL code is an inserted .\compile\programmable_prescalar_waveform.vhs
	--User can modify it ....

STIMULUS: process
begin  -- of stimulus process
--wait for <time to next event>; -- <current time>

	cs <= "000";
	clear <= '0';
	clk <= '0';
    wait for 50 ns; --0 fs
	clk <= '1';
    wait for 50 ns; --50 ns
	clk <= '0';
    wait for 50 ns; --100 ns
	clear <= '1';
	clk <= '1';
    wait for 50 ns; --150 ns
	clk <= '0';
    wait for 50 ns; --200 ns
	clk <= '1';
    wait for 50 ns; --250 ns
	clk <= '0';
    wait for 50 ns; --300 ns
	clk <= '1';
    wait for 50 ns; --350 ns
	clk <= '0';
    wait for 50 ns; --400 ns
	clk <= '1';
    wait for 50 ns; --450 ns
	cs <= "001";
	clk <= '0';
    wait for 50 ns; --500 ns
	clk <= '1';
    wait for 50 ns; --550 ns
	clk <= '0';
    wait for 50 ns; --600 ns
	clk <= '1';
    wait for 50 ns; --650 ns
	clk <= '0';
    wait for 50 ns; --700 ns
	clk <= '1';
    wait for 50 ns; --750 ns
	clk <= '0';
    wait for 50 ns; --800 ns
	clk <= '1';
    wait for 50 ns; --850 ns
	clk <= '0';
    wait for 50 ns; --900 ns
	clk <= '1';
    wait for 50 ns; --950 ns
	cs <= "010";
	clk <= '0';
    wait for 50 ns; --1 us
	clk <= '1';
    wait for 50 ns; --1050 ns
	clk <= '0';
    wait for 50 ns; --1100 ns
	clk <= '1';
    wait for 50 ns; --1150 ns
	clk <= '0';
    wait for 50 ns; --1200 ns
	clk <= '1';
    wait for 50 ns; --1250 ns
	clk <= '0';
    wait for 50 ns; --1300 ns
	clk <= '1';
    wait for 50 ns; --1350 ns
	clk <= '0';
    wait for 50 ns; --1400 ns
	clk <= '1';
    wait for 50 ns; --1450 ns
	cs <= "011";
	clk <= '0';
    wait for 50 ns; --1500 ns
	clk <= '1';
    wait for 50 ns; --1550 ns
	clk <= '0';
    wait for 50 ns; --1600 ns
	clk <= '1';
    wait for 50 ns; --1650 ns
	clk <= '0';
    wait for 50 ns; --1700 ns
	clk <= '1';
    wait for 50 ns; --1750 ns
	clk <= '0';
    wait for 50 ns; --1800 ns
	clk <= '1';
    wait for 50 ns; --1850 ns
	clk <= '0';
    wait for 50 ns; --1900 ns
	clk <= '1';
    wait for 50 ns; --1950 ns
	cs <= "100";
	clk <= '0';
    wait for 50 ns; --2 us
	clk <= '1';
    wait for 50 ns; --2050 ns
	clk <= '0';
    wait for 50 ns; --2100 ns
	clk <= '1';
    wait for 50 ns; --2150 ns
	clk <= '0';
    wait for 50 ns; --2200 ns
	clk <= '1';
    wait for 50 ns; --2250 ns
	clk <= '0';
    wait for 50 ns; --2300 ns
	clk <= '1';
    wait for 50 ns; --2350 ns
	clk <= '0';
    wait for 50 ns; --2400 ns
	clk <= '1';
    wait for 50 ns; --2450 ns
	cs <= "101";
	clk <= '0';
    wait for 50 ns; --2500 ns
	clk <= '1';
    wait for 50 ns; --2550 ns
	clk <= '0';
    wait for 50 ns; --2600 ns
	clk <= '1';
    wait for 50 ns; --2650 ns
	clk <= '0';
    wait for 50 ns; --2700 ns
	clk <= '1';
    wait for 50 ns; --2750 ns
	clk <= '0';
    wait for 50 ns; --2800 ns
	clk <= '1';
    wait for 50 ns; --2850 ns
	clk <= '0';
    wait for 50 ns; --2900 ns
	clk <= '1';
    wait for 50 ns; --2950 ns
	cs <= "110";
	clk <= '0';
--	end of stimulus events
	wait;
end process; -- end of stimulus process
	



	-- Add your stimulus here ...

end testbench;

configuration TESTBENCH_FOR_programmable_prescalar of programmable_prescalar_tb is
	for testbench
		for UUT : programmable_prescalar
			use entity work.programmable_prescalar(NetList);
		end for;
	end for;
end TESTBENCH_FOR_programmable_prescalar;

