configuration TIMING_FOR_decoder_3to8 of decoder_3to8_tb is
	for testbench
		for UUT : decoder_3to8
--
-- The user should replace : 
-- ENTITY_NAME with an	entity name from a backannotated VHDL file,
-- ARCH_NAME   with an architecture name from a backannotated VHDL file,
-- and uncomment the line below
--			use entity work.ENTITY_NAME (ARCH_NAME);
		end for;
	end for;
end TIMING_FOR_decoder_3to8;

